// // INSA : circular buffer used to store the first and last 
// module circular_buffer_om
// #(
//     parameter SIZE_BUFFER 10,
//     parameter SIZE_WORD 32
// )
// (
//     input logic       en_write,
//     input logic[31:0] find_in,
//     input logic[31:0] data_in,
//     output logic      data_in_memory
// );
//     data_in_memory
// endmodule
